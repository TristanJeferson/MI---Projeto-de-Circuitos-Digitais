module DecodificadorDisplay(bits, cadeia);

	input [3:0] bits;
	output reg [27:0] cadeia;
	
	always @(bits) begin
		case(bits)
			4'b0000: cadeia = 28'b0110000010010000110001111111;
			4'b0001:	cadeia = 28'b0110001011000011111111111111;
			4'b0010:	cadeia = 28'b0110001111000111111111111111;
			4'b0011: cadeia = 28'b0110001011000111111111111111;
			4'b0100: cadeia = 28'b0110001000100011111111111111;
			4'b0101: cadeia = 28'b0100100000100011111111111111;
			4'b0110: cadeia = 28'b0100100011000111111111111111;
			4'b0111: cadeia = 28'b0111000011000111111111111111;
			4'b1000: cadeia = 28'b1111111111111111111110000001;
			4'b1001: cadeia = 28'b1111111111111111111110010010;
			4'b1010: cadeia = 28'b1111111111111111111111001100;
			4'b1011: cadeia = 28'b1111111111111111111110100100;
			4'b1100: cadeia = 28'b1111111111111111111110100000;
			4'b1101: cadeia = 28'b1111111111111111111110000000;
			4'b1110: cadeia = 28'b0011000000100001000010000001;
			4'b1111: cadeia = 28'b1111111111111111111111111111;
		endcase
	end
endmodule