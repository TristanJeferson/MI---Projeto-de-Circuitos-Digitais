module main(CH7, CH6, CH5, CH4, CH3, CH2, CH1, B3, B0, CLK, RGB, BITS_DIGITOS, BITS_SEGMENTOS, LEDS);
	
	input CH7, CH6, CH5, CH4, CH3, CH2, CH1, B3, B0, CLK;
	
	
	wire CLK760HZ, CLK8S, CLK2S, CONFIRMA, INSERIR_CEDULA, LED1, LED2, LED3, LED4, LED5, LED6, LED7, LED8, LED9, LED10;
	wire [1:0] S_SENSORES, S_PAGAMENTO, S_ESCOLHA;
	wire [2:0] S_MAQUINA;
	wire [3:0] BITS_DISPLAY;
	wire [6:0] SAIDA_D_MAQUINA, SAIDA_D_SENSORES, SAIDA_D_PAGAMENTO, SAIDA_D_ESCOLHA;
	
	output [2:0] RGB;
	output [4:0] BITS_DIGITOS;
	output [6:0] BITS_SEGMENTOS;
	output [9:0] LEDS;
	
	
	DivisorFrequencia(CLK, CLK760HZ, CLK8S, CLK2S);
	LevelToPulse(B3, CLK760HZ, CONFIRMA);
	LevelToPulse(B0, CLK760HZ, INSERIR_CEDULA);
	MEFCafe(CLK760HZ, CONFIRMA, CLK8S, CLK2S, S_SENSORES, S_PAGAMENTO, S_ESCOLHA, SAIDA_D_MAQUINA, S_MAQUINA);
	MaquinaSensores(CLK760HZ, CLK8S, CH5, CH4, CH3, S_SENSORES, SAIDA_D_SENSORES);
	MaquinaPagamento(INSERIR_CEDULA, CLK8S, {CH7, CH6}, {CH2, CH1}, SAIDA_D_PAGAMENTO, S_PAGAMENTO);
	MaquinaEscolha(CLK760HZ, CLK8S, CONFIRMA, CH7, CH6, SAIDA_D_ESCOLHA, S_ESCOLHA);
	MuxSaidas(SAIDA_D_PAGAMENTO, SAIDA_D_SENSORES, SAIDA_D_ESCOLHA, SAIDA_D_MAQUINA, S_MAQUINA, BITS_DISPLAY);
	display(CLK760HZ, BITS_DISPLAY, BITS_DIGITOS, BITS_SEGMENTOS);
	
//	assign LED1 = (((!S_MAQUINA[2] && !S_MAQUINA[1]) || (S_MAQUINA[2] && S_MAQUINA[1])) && S_MAQUINA[0]);
//	assign LED2 = LED1;
//	assign LED3 = (((!S_MAQUINA[2] && !S_MAQUINA[0]) || (S_MAQUINA[2] && S_MAQUINA[0])) && S_MAQUINA[1]);
//	assign LED4 = LED3;
//	assign LED5 = (S_MAQUINA[1] && S_MAQUINA[0]);
//	assign LED6 = LED5;
//	assign LED7 = (S_MAQUINA[2] && S_MAQUINA[0]);
//	assign LED8 = LED7;
//	assign LED9 = (S_MAQUINA[2] && S_MAQUINA[1]);
//	assign LED10 = LED9;
	
	assign LEDS = {(((!S_MAQUINA[2] && !S_MAQUINA[1]) || (S_MAQUINA[2] && S_MAQUINA[1])) && S_MAQUINA[0]),
			(((!S_MAQUINA[2] && !S_MAQUINA[1]) || (S_MAQUINA[2] && S_MAQUINA[1])) && S_MAQUINA[0]),
			(((!S_MAQUINA[2] && !S_MAQUINA[0]) || (S_MAQUINA[2] && S_MAQUINA[0])) && S_MAQUINA[1]),
			(((!S_MAQUINA[2] && !S_MAQUINA[0]) || (S_MAQUINA[2] && S_MAQUINA[0])) && S_MAQUINA[1]),
			(S_MAQUINA[1] && S_MAQUINA[0]),
			(S_MAQUINA[1] && S_MAQUINA[0]),
			(S_MAQUINA[2] && S_MAQUINA[0]),
			(S_MAQUINA[2] && S_MAQUINA[0]),
			(S_MAQUINA[2] && S_MAQUINA[1]),
			(S_MAQUINA[2] && S_MAQUINA[1])};
	
	assign RGB = {(S_MAQUINA[2] && !S_MAQUINA[1]) || (!S_MAQUINA[2] && S_MAQUINA[0]) || (S_MAQUINA[1] && !S_MAQUINA[0]),
	(S_MAQUINA[1] || (!S_MAQUINA[1] && S_MAQUINA[0])),
	(!S_MAQUINA[2] && !S_MAQUINA[1] && !S_MAQUINA[0]) || (S_MAQUINA[2] && ((!S_MAQUINA[1] && S_MAQUINA[0]) || (S_MAQUINA[1] && !S_MAQUINA[0])))};


endmodule